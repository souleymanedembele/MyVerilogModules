/**
 * File              : RX.sv
 * Author            : Souleymane Dembele <sdembele@uw.edu>
 * Date              : 06.18.2023
 * Last Modified Date: 06.18.2023
 * Last Modified By  : Souleymane Dembele <sdembele@uw.edu>
 */
// this is the UART RX module
module RX (
    Clock,
    ClearN
);
endmodule
